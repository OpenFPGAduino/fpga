module matrix(
output AX_step_motor_0,
output AY_step_motor_0,
output BX_step_motor_0,
output BY_step_motor_0,
output AE_step_motor_0,
output BE_step_motor_0,

output AX_step_motor_1,
output AY_step_motor_1,
output BX_step_motor_1,
output BY_step_motor_1,
output AE_step_motor_1,
output BE_step_motor_1,

output AX_step_motor_2,
output AY_step_motor_2,
output BX_step_motor_2,
output BY_step_motor_2,
output AE_step_motor_2,
output BE_step_motor_2,

output AX_step_motor_3,
output AY_step_motor_3,
output BX_step_motor_3,
output BY_step_motor_3,
output AE_step_motor_3,
output BE_step_motor_3,

output HX_brush_motor_0,
output HY_brush_motor_0,

output HX_brush_motor_1,
output HY_brush_motor_1,

output HX_brush_motor_2,
output HY_brush_motor_2,

output HX_brush_motor_3,
output HY_brush_motor_3,

output sck_sht1x_sensor_0,
input dir_sht1x_sensor_0,
inout sda_sht1x_sensor_0,

inout PIN_0_PIOIN26_A,
inout PIN_1_PIOIN26_A,
inout PIN_2_PIOIN26_A,
inout PIN_3_PIOIN26_A,
inout PIN_4_PIOIN26_A,
inout PIN_5_PIOIN26_A,
inout PIN_6_PIOIN26_A,
inout PIN_7_PIOIN26_A,
inout PIN_8_PIOIN26_A,
inout PIN_9_PIOIN26_A,
inout PIN_10_PIOIN26_A,
inout PIN_11_PIOIN26_A,
inout PIN_12_PIOIN26_A,
inout PIN_13_PIOIN26_A,
inout PIN_14_PIOIN26_A,
inout PIN_15_PIOIN26_A,
inout PIN_16_PIOIN26_A,
inout PIN_17_PIOIN26_A,
inout PIN_18_PIOIN26_A,
inout PIN_19_PIOIN26_A,
inout PIN_20_PIOIN26_A,
inout PIN_21_PIOIN26_A,
inout PIN_22_PIOIN26_A,
inout PIN_23_PIOIN26_A,
inout PIN_24_PIOIN26_A,
inout PIN_25_PIOIN26_A,

inout PIN_0_PIOIN26_B,
inout PIN_1_PIOIN26_B,
inout PIN_2_PIOIN26_B,
inout PIN_3_PIOIN26_B,
inout PIN_4_PIOIN26_B,
inout PIN_5_PIOIN26_B,
inout PIN_6_PIOIN26_B,
inout PIN_7_PIOIN26_B,
inout PIN_8_PIOIN26_B,
inout PIN_9_PIOIN26_B,
inout PIN_10_PIOIN26_B,
inout PIN_11_PIOIN26_B,
inout PIN_12_PIOIN26_B,
inout PIN_13_PIOIN26_B,
inout PIN_14_PIOIN26_B,
inout PIN_15_PIOIN26_B,
inout PIN_16_PIOIN26_B,
inout PIN_17_PIOIN26_B,
inout PIN_18_PIOIN26_B,
inout PIN_19_PIOIN26_B,
inout PIN_20_PIOIN26_B,
inout PIN_21_PIOIN26_B,
inout PIN_22_PIOIN26_B,
inout PIN_23_PIOIN26_B,
inout PIN_24_PIOIN26_B,
inout PIN_25_PIOIN26_B,

inout PIN_0_PIO26_A,
inout PIN_1_PIO26_A,
inout PIN_2_PIO26_A,
inout PIN_3_PIO26_A,
inout PIN_4_PIO26_A,
inout PIN_5_PIO26_A,
inout PIN_6_PIO26_A,
inout PIN_7_PIO26_A,
inout PIN_8_PIO26_A,
inout PIN_9_PIO26_A,
inout PIN_10_PIO26_A,
inout PIN_11_PIO26_A,
inout PIN_12_PIO26_A,
inout PIN_13_PIO26_A,
inout PIN_14_PIO26_A,
inout PIN_15_PIO26_A,
inout PIN_16_PIO26_A,
inout PIN_17_PIO26_A,
inout PIN_18_PIO26_A,
inout PIN_19_PIO26_A,
inout PIN_20_PIO26_A,
inout PIN_21_PIO26_A,
inout PIN_22_PIO26_A,
inout PIN_23_PIO26_A,
inout PIN_24_PIO26_A,
inout PIN_25_PIO26_A,

inout PIN_0_PIO26_B,
inout PIN_1_PIO26_B,
inout PIN_2_PIO26_B,
inout PIN_3_PIO26_B,
inout PIN_4_PIO26_B,
inout PIN_5_PIO26_B,
inout PIN_6_PIO26_B,
inout PIN_7_PIO26_B,
inout PIN_8_PIO26_B,
inout PIN_9_PIO26_B,
inout PIN_10_PIO26_B,
inout PIN_11_PIO26_B,
inout PIN_12_PIO26_B,
inout PIN_13_PIO26_B,
inout PIN_14_PIO26_B,
inout PIN_15_PIO26_B,
inout PIN_16_PIO26_B,
inout PIN_17_PIO26_B,
inout PIN_18_PIO26_B,
inout PIN_19_PIO26_B,
inout PIN_20_PIO26_B,
inout PIN_21_PIO26_B,
inout PIN_22_PIO26_B,
inout PIN_23_PIO26_B,
inout PIN_24_PIO26_B,
inout PIN_25_PIO26_B,

input clock);
assign PIN_6_PIO26_A = AX_step_motor_1;
assign PIN_8_PIO26_A = AY_step_motor_1;
assign PIN_7_PIO26_A = BX_step_motor_1;
assign PIN_9_PIO26_A = BY_step_motor_1;
assign PIN_10_PIO26_A = AE_step_motor_1;
assign PIN_11_PIO26_A = BE_step_motor_1;
assign PIN_12_PIO26_A = AX_step_motor_2;
assign PIN_14_PIO26_A = AY_step_motor_2;
assign PIN_13_PIO26_A = BX_step_motor_2;
assign PIN_15_PIO26_A = BY_step_motor_2;
assign PIN_16_PIO26_A = AE_step_motor_2;
assign PIN_17_PIO26_A = BE_step_motor_2;
assign PIN_0_PIO26_B = HX_brush_motor_0;
assign PIN_1_PIO26_B = HY_brush_motor_0;
endmodule
